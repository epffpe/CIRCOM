S 1 3
.lib cmos6tm.mod

.param ancho=10u
.param largo=10u

.param amp=50m
.param frec=1k
M1 vdd G vss vss modn w={ancho} l={largo}

VSS vss 0 0 DC 0

VDD vdd vss  5 DC 5
Vbias pol vss  3 DC 3
Vin G pol sin(0 {amp} {frec})
.op
.tran 0 5m 0.01m

.probe

.end
