E 1_44
.lib cmos6tm.mod
.param ancho=150u
.param largo=0.35u
M1		D	G	0	0	modn	 w={ancho} 	l={largo} ; transistor principal

Rl		vcc	D	1k
Cl		vcc	D	7.78p
Ll		D2		D	1nH
Cs		vcc	D2	10u
Vcc	vcc	0	5V
Vbias	g1		0	1.08V
Vin	G		g1	DC 0	AC 100m	SIN(0 100m 1G)

.op
.tran 0.1n 100n
*.ac DEC 5k	1Meg	7G
.probe
.end
