S 1 2
.lib cmos6tm.mod

.param ancho=10u
.param largo=10u

M1 vdd G vss vss modn w={ancho} l={largo}

VSS vss 0 0 DC 0

VDD vdd vss  5 DC 5
Vbias G vss  1 DC 1

.dc Vbias 0 5 0.5

.probe

.end
