S 2 17
.lib cmos6tm.mod

.param ancho=150u
.param largo=0.35u

.param amp=4
.param amp2=2
.param f1=1Meg
.param f2=1.8Meg
.param fas1=0
.param fas2=90
M1 vdd G out vss modn w={ancho} l={largo}



ibias out vss sin(1m 0.5m {f1})

VSS vss 0 0 DC 0
VDD vdd vss  5 DC 5
Vbias G vss  2.5 DC 2.5

.op
.tran 0 5u 0.01u
.probe

.end
