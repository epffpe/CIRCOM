S 1 4
.lib cmos6tm.mod

.param ancho=10u
.param largo=10u

.param amp=4
.param frec=1k
M1 vdd G vss vss modn w={ancho} l={largo}

VSS vss 0 0 DC 0

VDD vdd vss  5 DC 5
Vbias pol vss  3 DC 3
Vin G pol sin(0 {amp} {frec})
.op
.tran 0 12m 0.05m

.probe

.end
