S 2 16
.lib cmos6tm.mod

.param ancho=150u
.param largo=0.35u

.param amp=4
.param amp2=2
.param f1=1Meg
.param f2=1.8Meg
.param fas1=0
.param fas2=90
M1 vdd G out vss modn w={ancho} l={largo}




Ibias out vss 1m DC 1m
VSS vss 0 0 DC 0
VDD vdd vss  5 DC 5
Vbias pol vss  2.5 DC 2.5
vgsignal1 pol in2 sin(0 {amp} {f1} 0 0 {fas1})
vgsignal2 in2 G sin(0 {amp2} {f2} 0 0 {fas2})
.op
.tran 0 5u 0.01u
.probe

.end
