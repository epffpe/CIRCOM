S 2 13
.lib cmos6tm.mod

.param ancho=150u
.param largo=0.35u

.param ampl=4
.param freq=1k
M1 out G vss vss modn w={ancho} l={largo}
Rl vdd out 1k
VSS vss 0 0 DC 0

VDD vdd vss  5 DC 5
Vbias pol vss  1.08 DC 1.08
Vin pol G sin(0 {ampl} {freq}) AC 0.05
.op
.ac dec 100 10 1000G

.probe

.end
